module fht_but #(parameter D_BIT = 17, W_BIT = 12)(
	input iCLK,
	input iRESET,
	
//	input iSEL,
	
	input signed [D_BIT - 1 : 0] iX_0,
	input signed [D_BIT - 1 : 0] iX_1,
	input signed [D_BIT - 1 : 0] iX_2,
	
	input signed [W_BIT - 1 : 0] iSIN,
	input signed [W_BIT - 1 : 0] iCOS,
	
	output signed [D_BIT - 1 : 0] oY_0,
	output signed [D_BIT - 1 : 0] oY_1
);

reg signed [D_BIT - 1 : 0] sum_mul;

reg signed [D_BIT - 1 : 0] sum_buf;
reg signed [D_BIT - 1 : 0] sub_buf;

wire signed [D_BIT + W_BIT : 0] EXT_SUM_MUL = iX_1 * iCOS + iX_2 * iSIN + 2'sd1;

//wire signed [D_BIT - 1 : 0] MUX_SUM = iSEL ? (iX_1) : (mul_cos_buf + mul_sin_buf); // for '0' stage
//wire signed [D_BIT - 1 : 0] MUX_SUB = iSEL ? (iX_1) : (mul_cos_buf - mul_sin_buf);

wire signed [D_BIT : 0] EXT_SUM = iX_0 + sum_mul + 2'sd1;
wire signed [D_BIT : 0] EXT_SUB = iX_0 - sum_mul + 2'sd1;

always@(posedge iCLK or negedge iRESET)begin
	if(!iRESET) sum_mul <= 0;
	else sum_mul <= EXT_SUM_MUL[D_BIT + W_BIT - 2 : W_BIT - 1];
end

always@(posedge iCLK or negedge iRESET)begin
	if(!iRESET)
		begin
			sum_buf <= 0;
			sub_buf <= 0;
		end
	else
		begin
			sum_buf <= EXT_SUM[D_BIT : 1];
			sub_buf <= EXT_SUB[D_BIT : 1];
		end
end

assign oY_0 = sum_buf;
assign oY_1 = sub_buf;

endmodule 
typedef integer unsigned	uint32_t;
typedef shortint unsigned	uint16_t;

typedef real		float64_t;
typedef shortreal	float32_t;


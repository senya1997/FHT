
`include "TransformRAM.svh"

function automatic void TransformRAM::Save_RAM_data(string name, bit ram_sel); // 0 - RAM(A), 1 - RAM(B)

endfunction
